module vpu_core(
  input wire clk,
  input wire rst,
  input [31:0] vram_addr,
  input [31:0] tileram_addr,
);

endmodule
