module board (
  input  wire        clk,
  input  wire        rst_n,

  input  wire        clk,
  input  wire        rst_n,
);

endmodule
