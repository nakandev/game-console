package gameconsole_pkg;

parameter SCREEN_W      = 320;
parameter SCREEN_H      = 240;
parameter SCREEN_HBLANK =  80;
parameter SCREEN_VBLANK =  80;
parameter SP_ADDR_W     =  10;
parameter SP_DATA_W     =  32;
parameter MAP_ADDR_W    =  11;
parameter MAP_DATA_W    =  16;
parameter TILE_ADDR_W   =  15;
parameter TILE_DATA_W   =   8;
parameter PAL_ADDR_W    =   8;
parameter PAL_DATA_W    =  32;

endpackage
